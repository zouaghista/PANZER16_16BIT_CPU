`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:33:17 06/30/2024 
// Design Name: 
// Module Name:    Mux16_4 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Mux16_4(
    input Sel,
    input [15:0] Input1,
    input [15:0] Input2,
    input [15:0] Input3,
    input [15:0] Input4,
    output [15:0] Output
    );


endmodule
