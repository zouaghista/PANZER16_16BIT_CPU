`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    03:51:06 06/02/2024 
// Design Name: 
// Module Name:    DeMux16_2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module DeMux16_2(
    input sel,
    output [15:0] output1,
    output [15:0] output2,
    input [15:0] Input
    );


endmodule
